package CustomReg;

typedef 640 MAX_CUSTOM_REG_SIZE;
Bit#(10) max_custom_reg_size = 640;

endpackage