package CustomReg;

typedef 64 MAX_CUSTOM_REG_SIZE;
Bit#(7) max_custom_reg_size = 64;

endpackage